`timescale 1ns/1ns

module AND(
		input A,B,
		output Sal
);

assign Sal = A & B;

endmodule 